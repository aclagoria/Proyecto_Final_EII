library IEEE;
use IEEE.std_logic_1164.all;
package pkg_tabla_caracteres is
    type Tabla_256x64 is array (0 to 256) of std_logic_vector (64 downto 0);
end package;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.pkg_tabla_caracteres.all;

entity tabla_caracteres is
    generic (
        constant fuente : tabla_fuente  := (others=>(others=>'0')));
    port(
        dir  : in std_logic_vector (7 downto 0);
        dato : out std_logic_vector (63 downto 0));
end tabla_caracteres;

architecture solucion of tabla_caracteres is
    constant fuente : tabla_fuente :=(
    0=> x"0000000000000000",
    1=> x"7e81a581bd99817e",
    2=> x"7effdbffc3e7ff7e",
    3=> x"6cfefefe7c381000",
    4=> x"10387cfe7c381000",
    5=> x"387c38fefed61038",
    6=> x"1010387cfe7c1038",
    7=> x"0000183c3c180000",
    8=> x"ffffe7c3c3e7ffff",
    9=> x"003c664242663c00",
    10=> x"ffc399bdbd99c3ff",
    11=> x"0f070f7dcccccc78",
    12=> x"3c6666663c187e18",
    13=> x"3f333f303070f0e0",
    14=> x"7f637f636367e6c0",
    15=> x"995a3ce7e73c5a99",
    16=> x"80e0f8fef8e08000",
    17=> x"020e3efe3e0e0200",
    18=> x"183c7e18187e3c18",
    19=> x"6666666666006600",
    20=> x"7fdbdb7b1b1b1b00",
    21=> x"7ec378cccc788cf8",
    22=> x"000000007e7e7e00",
    23=> x"183c7e187e3c18ff",
    24=> x"183c7e1818181800",
    25=> x"181818187e3c1800",
    26=> x"00180cfe0c180000",
    27=> x"003060fe60300000",
    28=> x"0000c0c0c0fe0000",
    29=> x"002466ff66240000",
    30=> x"00183c7effff0000",
    31=> x"00ffff7e3c180000",
    32=> x"0000000000000000",
    33=> x"3078783030003000",
    34=> x"6c6c6c0000000000",
    35=> x"6c6cfe6cfe6c6c00",
    36=> x"307cc0780cf83000",
    37=> x"00c6cc183066c600",
    38=> x"386c3876dccc7600",
    39=> x"6060c00000000000",
    40=> x"1830606060301800",
    41=> x"6030181818306000",
    42=> x"00663cff3c660000",
    43=> x"003030fc30300000",
    44=> x"0000000000703060",
    45=> x"000000fc00000000",
    46=> x"0000000000303000",
    47=> x"060c183060c08000",
    48=> x"78ccdcfceccc7800",
    49=> x"30f030303030fc00",
    50=> x"78cc0c3860ccfc00",
    51=> x"78cc0c380ccc7800",
    52=> x"1c3c6cccfe0c0c00",
    53=> x"fcc0f80c0ccc7800",
    54=> x"3860c0f8cccc7800",
    55=> x"fccc0c1830606000",
    56=> x"78cccc78cccc7800",
    57=> x"78cccc7c0c187000",
    58=> x"0000303000303000",
    59=> x"0000303000703060",
    60=> x"183060c060301800",
    61=> x"0000fc00fc000000",
    62=> x"6030180c18306000",
    63=> x"78cc0c1830003000",
    64=> x"7cc6dededec07800",
    65=> x"3078ccccfccccc00",
    66=> x"fc66667c6666fc00",
    67=> x"3c66c0c0c0663c00",
    68=> x"fc6c6666666cfc00",
    69=> x"fe6268786862fe00",
    70=> x"fe6268786860f000",
    71=> x"3c66c0c0ce663e00",
    72=> x"ccccccfccccccc00",
    73=> x"7830303030307800",
    74=> x"1e0c0c0ccccc7800",
    75=> x"e6666c786c66e600",
    76=> x"f06060606266fe00",
    77=> x"c6eefed6c6c6c600",
    78=> x"c6e6f6decec6c600",
    79=> x"386cc6c6c66c3800",
    80=> x"fc66667c6060f000",
    81=> x"78ccccccdc781c00",
    82=> x"fc66667c786ce600",
    83=> x"78cce0381ccc7800",
    84=> x"fcb4303030307800",
    85=> x"ccccccccccccfc00",
    86=> x"cccccccccc783000",
    87=> x"c6c6c6d6feeec600",
    88=> x"c6c66c386cc6c600",
    89=> x"cccccc7830307800",
    90=> x"fecc983062c6fe00",
    91=> x"7860606060607800",
    92=> x"c06030180c060200",
    93=> x"7818181818187800",
    94=> x"10386cc600000000",
    95=> x"00000000000000ff",
    96=> x"3030180000000000",
    97=> x"0000780c7ccc7600",
    98=> x"e0607c666666bc00",
    99=> x"000078ccc0cc7800",
    100=> x"1c0c0c7ccccc7600",
    101=> x"000078ccfcc07800",
    102=> x"386c60f06060f000",
    103=> x"000076cccc7c0cf8",
    104=> x"e0606c766666e600",
    105=> x"3000703030307800",
    106=> x"180078181818d870",
    107=> x"e060666c786ce600",
    108=> x"7030303030307800",
    109=> x"0000ecfed6c6c600",
    110=> x"0000f8cccccccc00",
    111=> x"000078cccccc7800",
    112=> x"0000dc66667c60f0",
    113=> x"000076cccc7c0c1e",
    114=> x"0000d86c6c60f000",
    115=> x"00007cc0780cf800",
    116=> x"10307c3030341800",
    117=> x"0000cccccccc7600",
    118=> x"0000cccccc783000",
    119=> x"0000c6c6d6fe6c00",
    120=> x"0000c66c386cc600",
    121=> x"0000cccccc7c0cf8",
    122=> x"0000fc983064fc00",
    123=> x"1c3030e030301c00",
    124=> x"1818180018181800",
    125=> x"e030301c3030e000",
    126=> x"76dc000000000000",
    127=> x"10386cc6c6c6fe00",
    128=> x"78ccc0cc78180c78",
    129=> x"00cc00cccccc7e00",
    130=> x"1c0078ccfcc07800",
    131=> x"7ec33c063e663f00",
    132=> x"cc00780c7ccc7e00",
    133=> x"e000780c7ccc7e00",
    134=> x"3030780c7ccc7e00",
    135=> x"00007cc0c07c063c",
    136=> x"7ec33c667e603c00",
    137=> x"cc0078ccfcc07800",
    138=> x"e00078ccfcc07800",
    139=> x"cc00703030307800",
    140=> x"7cc6381818183c00",
    141=> x"e000703030307800",
    142=> x"cc3078ccccfccc00",
    143=> x"30300078ccfccc00",
    144=> x"1c00fc607860fc00",
    145=> x"00007f0c7fcc7f00",
    146=> x"3e6cccfeccccce00",
    147=> x"78cc0078cccc7800",
    148=> x"00cc0078cccc7800",
    149=> x"00e00078cccc7800",
    150=> x"78cc00cccccc7e00",
    151=> x"00e000cccccc7e00",
    152=> x"00cc00ccccfc0cf8",
    153=> x"c6387cc6c67c3800",
    154=> x"cc00cccccccc7800",
    155=> x"18187ec0c07e1818",
    156=> x"386c64f060e6fc00",
    157=> x"cccc78fc30fc3000",
    158=> x"f0d8d8f4ccdecc0e",
    159=> x"0e1b187e1818d870",
    160=> x"1c00780c7ccc7e00",
    161=> x"3800703030307800",
    162=> x"001c0078cccc7800",
    163=> x"001c00cccccc7e00",
    164=> x"00f800f8cccccc00",
    165=> x"fc00ccecfcdccc00",
    166=> x"3c6c6c3e007e0000",
    167=> x"3c66663c007e0000",
    168=> x"30003060c0cc7800",
    169=> x"000000fcc0c00000",
    170=> x"000000fc0c0c0000",
    171=> x"c6ccd83e63ce981f",
    172=> x"c6ccd8f367cf9f03",
    173=> x"00180018183c3c18",
    174=> x"003366cc66330000",
    175=> x"00cc663366cc0000",
    176=> x"2288228822882288",
    177=> x"55aa55aa55aa55aa",
    178=> x"dd77dd77dd77dd77",
    179=> x"1818181818181818",
    180=> x"18181818f8181818",
    181=> x"1818f818f8181818",
    182=> x"36363636f6363636",
    183=> x"00000000fe363636",
    184=> x"0000f818f8181818",
    185=> x"3636f606f6363636",
    186=> x"3636363636363636",
    187=> x"0000fe06f6363636",
    188=> x"3636f606fe000000",
    189=> x"36363636fe000000",
    190=> x"1818f818f8000000",
    191=> x"00000000f8181818",
    192=> x"181818181f000000",
    193=> x"18181818ff000000",
    194=> x"00000000ff181818",
    195=> x"181818181f181818",
    196=> x"00000000ff000000",
    197=> x"18181818ff181818",
    198=> x"18181f181f181818",
    199=> x"3636363637363636",
    200=> x"363637303f000000",
    201=> x"00003f3037363636",
    202=> x"3636f700ff000000",
    203=> x"0000ff00f7363636",
    204=> x"3636373037363636",
    205=> x"0000ff00ff000000",
    206=> x"3636f700f7363636",
    207=> x"1818ff00ff000000",
    208=> x"36363636ff000000",
    209=> x"0000ff00ff181818",
    210=> x"00000000ff363636",
    211=> x"363636363f000000",
    212=> x"18181f181f000000",
    213=> x"00001f181f181818",
    214=> x"000000003f363636",
    215=> x"36363636f7363636",
    216=> x"1818ff00ff181818",
    217=> x"18181818f8000000",
    218=> x"000000001f181818",
    219=> x"ffffffffffffffff",
    220=> x"00000000ffffffff",
    221=> x"f0f0f0f0f0f0f0f0",
    222=> x"0f0f0f0f0f0f0f0f",
    223=> x"ffffffff00000000",
    224=> x"000076dcc8dc7600",
    225=> x"0078ccf8ccf8c0c0",
    226=> x"00fec6c0c0c0c000",
    227=> x"00fe6c6c6c6c6c00",
    228=> x"fe6630183066fe00",
    229=> x"00007ecccccc7800",
    230=> x"00666666667c60c0",
    231=> x"0076dc1818181800",
    232=> x"fc3078cccc7830fc",
    233=> x"386cc6fec66c3800",
    234=> x"386cc6c66c6cee00",
    235=> x"1c30187ccccc7800",
    236=> x"00007edbdb7e0000",
    237=> x"060c7edbdb7e60c0",
    238=> x"3c60c0fcc0603c00",
    239=> x"78cccccccccccc00",
    240=> x"00fc00fc00fc0000",
    241=> x"3030fc303000fc00",
    242=> x"603018306000fc00",
    243=> x"183060301800fc00",
    244=> x"0e1b1b1818181818",
    245=> x"1818181818d8d870",
    246=> x"303000fc00303000",
    247=> x"00729c00729c0000",
    248=> x"386c6c3800000000",
    249=> x"0000001818000000",
    250=> x"0000000018000000",
    251=> x"0f0c0c0cec6c3c1c",
    252=> x"786c6c6c6c000000",
    253=> x"780c38607c000000",
    254=> x"00003c3c3c3c0000",
    255=> x"0000000000000000");
begin

dato <= fuente(to_integer(dir)); 

end solucion;
